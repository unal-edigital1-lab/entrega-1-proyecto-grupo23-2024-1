
module sensor(
  
  
  
  
  
  );




  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
endmodule